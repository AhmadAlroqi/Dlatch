`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/18/2024 02:37:39 PM
// Design Name: 
// Module Name: mux
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux #(parameter n=4 )(

input logic [n-1:0]x,
input logic [n-1:0]y,
input logic s,
output logic [n-1:0]z

    );
    
always @ (*)
begin 
 if (s==0)
         z=x;
 else 
         z=y;
    
   end  
   
endmodule
